module main

fn add(a, b mut int) int {
    c := a + b
}

fn main() {
    print(a)
}
