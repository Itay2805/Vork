module main

const Pi = 3.14

fn main() {
    assert Pi == 3.14
}
