module time
