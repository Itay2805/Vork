module main

fn main() {
    mut arr := [1,2,3,4]
    arr[0] = 12
    print(arr[0])
}
