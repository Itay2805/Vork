module main

fn test(arr []int) {
    print(arr.len)
}

fn main() {
    test([[1,2,3].len]int)
}
