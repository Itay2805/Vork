module main

fn add(a, b int) int {
    return a + b
}

fn main() {
    a := add(1, 2)
    print(a)
}
