module main

import bitfield
import rand

fn main() {
}
