module main

fn add(a, b int) int {
    c := a + b
    return c
}

fn main() {
    c := add(12, 12)
    print(c)
}
