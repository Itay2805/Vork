module time

fn C.ticks() i64
pub fn ticks() i64 {
    return C.ticks()
}
