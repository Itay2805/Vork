module main

import bitfield
import rand
import time

fn main() {
}
