module main

import bitfield

fn main() {
    mut bf := bitfield.new(32)
    print(bf.getbit(0))
}
