module main

import bitfield

fn main() {
}
